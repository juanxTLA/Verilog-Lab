`timescale 1ns/1ps
module tb_SearchTable();
    reg           reset;
    reg            req;
    reg [47:0]    search;
    reg            opReq;
    reg [1:0]     opCode;
    reg [47:0]    opSearch;
    reg [15:0]    opResult;
    reg            clk;
    wire           opRdy;
    wire           rdy;
    wire           found;
    wire           done;
    wire [15:0]    result;
    wire           opErr;
    wire [10:0]    numEntries;

    initial begin
        opSearch = 48'h96;
        opReq    = 1'b1;
        opResult = 16'd68;
        clk = 0;
        opCode = 2'b00;
        req = 0;
        search = 48'h84;
    end


    always #5  clk = ~clk;
    always begin
        
        #20; opSearch = 48'h84; opResult = 16'd1;
        #20; opSearch = 48'h97; opResult = 16'd2;
        #20; opSearch = 48'h57; opResult = 16'd3;
        #20; opSearch = 48'h1; opResult = 16'd4;
        #20; opCode = 2'b01; opSearch = 48'h57;
        #20; opCode = 2'b10; opResult = 16'h89; opSearch = 48'h1;
        #20; opReq = 0; req = 1;
        #20; opReq = 1; req = 0; opCode = 2'b11; 

    end

    SearchTable uut(
        reset,
        req,
        search,
        opReq,
        opCode,
        opSearch,
        opResult,
        clk,
        opRdy,
        rdy,
        found,
        done,
        result,
        opErr,
        numEntries
    );
endmodule